LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Parallel4BitDecoder IS
  PORT (x: IN STD_LOGIC_VECTOR(7 downto 0);
        m:   OUT STD_LOGIC_VECTOR(3 downto 0));
END Parallel4BitDecoder;

ARCHITECTURE structure OF Parallel4BitDecoder IS

BEGIN
  

END structure;

ENTITY 

